typedef uvm_sequencer#(write_tx) write_sqr;
